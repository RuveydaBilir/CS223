`timescale 1ns / 1ps
module TB_Mux4to1;
reg d0, d1, d2, d3, s0, s1;
wire y;

Mux4to1 dut(.d0(d0), .d1(d1), .d2(d2), .d3(d3), .s0(s0), .s1(s1), .y(y) );

initial begin
 #100; d0 = 0; d1 = 0; d2 = 0; d3 = 0; s0 = 0; s1 = 0;
 #100; d0 = 0; d1 = 0; d2 = 0; d3 = 0; s0 = 0; s1 = 1;
 #100; d0 = 0; d1 = 0; d2 = 0; d3 = 0; s0 = 1; s1 = 0;
 #100; d0 = 0; d1 = 0; d2 = 0; d3 = 0; s0 = 1; s1 = 1;
 #100; d0 = 0; d1 = 0; d2 = 0; d3 = 1; s0 = 0; s1 = 0;
 #100; d0 = 0; d1 = 0; d2 = 0; d3 = 1; s0 = 0; s1 = 1;
 #100; d0 = 0; d1 = 0; d2 = 0; d3 = 1; s0 = 1; s1 = 0;
 #100; d0 = 0; d1 = 0; d2 = 0; d3 = 1; s0 = 1; s1 = 1;
 #100; d0 = 0; d1 = 0; d2 = 1; d3 = 0; s0 = 0; s1 = 0;
 #100; d0 = 0; d1 = 0; d2 = 1; d3 = 0; s0 = 0; s1 = 1;
 #100; d0 = 0; d1 = 0; d2 = 1; d3 = 0; s0 = 1; s1 = 0;
 #100; d0 = 0; d1 = 0; d2 = 1; d3 = 0; s0 = 1; s1 = 1;
 #100; d0 = 0; d1 = 0; d2 = 1; d3 = 1; s0 = 0; s1 = 0;
 #100; d0 = 0; d1 = 0; d2 = 1; d3 = 1; s0 = 0; s1 = 1;
 #100; d0 = 0; d1 = 0; d2 = 1; d3 = 1; s0 = 1; s1 = 0;
 #100; d0 = 0; d1 = 0; d2 = 1; d3 = 1; s0 = 1; s1 = 1;
 #100; d0 = 0; d1 = 1; d2 = 0; d3 = 0; s0 = 0; s1 = 0;
 #100; d0 = 0; d1 = 1; d2 = 0; d3 = 0; s0 = 0; s1 = 1;
 #100; d0 = 0; d1 = 1; d2 = 0; d3 = 0; s0 = 1; s1 = 0;
 #100; d0 = 0; d1 = 1; d2 = 0; d3 = 0; s0 = 1; s1 = 1;
 #100; d0 = 0; d1 = 1; d2 = 0; d3 = 1; s0 = 0; s1 = 0;
 #100; d0 = 0; d1 = 1; d2 = 0; d3 = 1; s0 = 0; s1 = 1;
 #100; d0 = 0; d1 = 1; d2 = 0; d3 = 1; s0 = 1; s1 = 0;
 #100; d0 = 0; d1 = 1; d2 = 0; d3 = 1; s0 = 1; s1 = 1;
 #100; d0 = 0; d1 = 1; d2 = 1; d3 = 0; s0 = 0; s1 = 0;
 #100; d0 = 0; d1 = 1; d2 = 1; d3 = 0; s0 = 0; s1 = 1;
 #100; d0 = 0; d1 = 1; d2 = 1; d3 = 0; s0 = 1; s1 = 0;
 #100; d0 = 0; d1 = 1; d2 = 1; d3 = 0; s0 = 1; s1 = 1;
 #100; d0 = 0; d1 = 1; d2 = 1; d3 = 1; s0 = 0; s1 = 0;
 #100; d0 = 0; d1 = 1; d2 = 1; d3 = 1; s0 = 0; s1 = 1;
 #100; d0 = 0; d1 = 1; d2 = 1; d3 = 1; s0 = 1; s1 = 0;
 #100; d0 = 0; d1 = 1; d2 = 1; d3 = 1; s0 = 1; s1 = 1;
 #100; d0 = 1; d1 = 0; d2 = 0; d3 = 0; s0 = 0; s1 = 0;
 #100; d0 = 1; d1 = 0; d2 = 0; d3 = 0; s0 = 0; s1 = 1;
 #100; d0 = 1; d1 = 0; d2 = 0; d3 = 0; s0 = 1; s1 = 0;
 #100; d0 = 1; d1 = 0; d2 = 0; d3 = 0; s0 = 1; s1 = 1;
 #100; d0 = 1; d1 = 0; d2 = 0; d3 = 1; s0 = 0; s1 = 0;
 #100; d0 = 1; d1 = 0; d2 = 0; d3 = 1; s0 = 0; s1 = 1;
 #100; d0 = 1; d1 = 0; d2 = 0; d3 = 1; s0 = 1; s1 = 0;
 #100; d0 = 1; d1 = 0; d2 = 0; d3 = 1; s0 = 1; s1 = 1;
 #100; d0 = 1; d1 = 0; d2 = 1; d3 = 0; s0 = 0; s1 = 0;
 #100; d0 = 1; d1 = 0; d2 = 1; d3 = 0; s0 = 0; s1 = 1;
 #100; d0 = 1; d1 = 0; d2 = 1; d3 = 0; s0 = 1; s1 = 0;
 #100; d0 = 1; d1 = 0; d2 = 1; d3 = 0; s0 = 1; s1 = 1;
 #100; d0 = 1; d1 = 0; d2 = 1; d3 = 1; s0 = 0; s1 = 0;
 #100; d0 = 1; d1 = 0; d2 = 1; d3 = 1; s0 = 0; s1 = 1;
 #100; d0 = 1; d1 = 0; d2 = 1; d3 = 1; s0 = 1; s1 = 0;
 #100; d0 = 1; d1 = 0; d2 = 1; d3 = 1; s0 = 1; s1 = 1;
 #100; d0 = 1; d1 = 1; d2 = 0; d3 = 0; s0 = 0; s1 = 0;
 #100; d0 = 1; d1 = 1; d2 = 0; d3 = 0; s0 = 0; s1 = 1;
 #100; d0 = 1; d1 = 1; d2 = 0; d3 = 0; s0 = 1; s1 = 0;
 #100; d0 = 1; d1 = 1; d2 = 0; d3 = 0; s0 = 1; s1 = 1;
 #100; d0 = 1; d1 = 1; d2 = 0; d3 = 1; s0 = 0; s1 = 0;
 #100; d0 = 1; d1 = 1; d2 = 0; d3 = 1; s0 = 0; s1 = 1;
 #100; d0 = 1; d1 = 1; d2 = 0; d3 = 1; s0 = 1; s1 = 0;
 #100; d0 = 1; d1 = 1; d2 = 0; d3 = 1; s0 = 1; s1 = 1;
 #100; d0 = 1; d1 = 1; d2 = 1; d3 = 0; s0 = 0; s1 = 0;
 #100; d0 = 1; d1 = 1; d2 = 1; d3 = 0; s0 = 0; s1 = 1;
 #100; d0 = 1; d1 = 1; d2 = 1; d3 = 0; s0 = 1; s1 = 0;
 #100; d0 = 1; d1 = 1; d2 = 1; d3 = 0; s0 = 1; s1 = 1;
 #100; d0 = 1; d1 = 1; d2 = 1; d3 = 1; s0 = 0; s1 = 0;
 #100; d0 = 1; d1 = 1; d2 = 1; d3 = 1; s0 = 0; s1 = 1;
 #100; d0 = 1; d1 = 1; d2 = 1; d3 = 1; s0 = 1; s1 = 0;
 #100; d0 = 1; d1 = 1; d2 = 1; d3 = 1; s0 = 1; s1 = 1;
end
endmodule
