`timescale 1ns / 1ps
module OneDisplay(
    input logic clk,
    input logic reset,
    input logic [3:0] number,
    output logic [6:0] seg
);
    
endmodule
