`timescale 1ns / 1ps
module TB_FunctionF;
    reg a,b,c,d,e;
    wire f;
FunctionF uut(.a(a), .b(b), .c(c), .d(d), .e(e), .f(f));

initial begin
#100 a=0; b=0; c=0; d=0; e=0;
#100 a=0; b=0; c=0; d=0; e=1;
#100 a=0; b=0; c=0; d=1; e=0;
#100 a=0; b=0; c=0; d=1; e=1;
#100 a=0; b=0; c=1; d=0; e=0;
#100 a=0; b=0; c=1; d=0; e=1;
#100 a=0; b=0; c=1; d=1; e=0;
#100 a=0; b=0; c=1; d=1; e=1;

#100 a=0; b=1; c=0; d=0; e=0;
#100 a=0; b=1; c=0; d=0; e=1;
#100 a=0; b=1; c=0; d=1; e=0;
#100 a=0; b=1; c=0; d=1; e=1;
#100 a=0; b=1; c=1; d=0; e=0;
#100 a=0; b=1; c=1; d=0; e=1;
#100 a=0; b=1; c=1; d=1; e=0;
#100 a=0; b=1; c=1; d=1; e=1;

#100 a=1; b=0; c=0; d=0; e=0;
#100 a=1; b=0; c=0; d=0; e=1;
#100 a=1; b=0; c=0; d=1; e=0;
#100 a=1; b=0; c=0; d=1; e=1;
#100 a=1; b=0; c=1; d=0; e=0;
#100 a=1; b=0; c=1; d=0; e=1;
#100 a=1; b=0; c=1; d=1; e=0;
#100 a=1; b=0; c=1; d=1; e=1;

#100 a=1; b=1; c=0; d=0; e=0;
#100 a=1; b=1; c=0; d=0; e=1;
#100 a=1; b=1; c=0; d=1; e=0;
#100 a=1; b=1; c=0; d=1; e=1;
#100 a=1; b=1; c=1; d=0; e=0;
#100 a=1; b=1; c=1; d=0; e=1;
#100 a=1; b=1; c=1; d=1; e=0;
#100 a=1; b=1; c=1; d=1; e=1;

end
endmodule
